module v1

pub struct PrevisaOceanica {
pub:
	cidade        string
	estado        string
	atualizado_em string
	ondas         []Ondas
}
