module v1

pub struct DadoOndas {
pub:
	vento              f32
	direcao_vento      string
	direcao_vento_desc string
	altura_onda        f32
	direcao_onda       string
	direcao_onda_desc  string
	agitacao           string
	hora               string
}
