module v1

pub struct Ddd {
pub:
	state  string
	cities []string
}
