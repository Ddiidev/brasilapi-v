module v1

pub enum TiposVeiculo {
	caminhoes
	carros
	motos
}
