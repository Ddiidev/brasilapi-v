module v1

pub struct Dimension {
pub:
	width f64
	height f64
	unit string
}
