module v1

pub struct Ondas {
pub:
	data        string
	dados_ondas []DadoOndas
}
