module errors

pub struct FeriadosNacionaisError {
	Error
	pub:
	message string
	@type   string
	name    string
}
