module v1

pub struct Cidade {
pub:
	nome   string
	estado string
	id     int
}
