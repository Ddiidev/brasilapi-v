module v1

pub struct Previsiao {
pub:
	cidade        string
	estado        string
	atualizado_em string
	clima         []Clima
}
