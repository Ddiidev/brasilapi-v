module v1

pub struct IBGE {
pub:
	nome        string
	codigo_ibge string
}
