module v1

pub struct Taxa {
pub:
	nome  string
	valor f32
}
