module v2

pub struct Coordinates {
pub:
	longitude string
	latitude  string
}
