module v1

// Classificação Nacional de Atividades Econômicas Secundárias da empresa.
pub struct CnaesSecundarios {
	pub:
	codigo    int
	descricao string
}
