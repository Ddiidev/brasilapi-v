module v1

pub struct DadoOndas {
pub:
	vento              float
	direcao_vento      string
	direcao_vento_desc string
	altura_onda        float
	direcao_onda       string
	direcao_onda_desc  string
	agitacao           string
	hora               string
}
