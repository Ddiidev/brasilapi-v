module v1

pub struct FipeMarcas {
pub:
	nome  string
	valor i64
}
