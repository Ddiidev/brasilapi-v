module v2

pub struct Cep {
pub:
	cep          string
	state        string
	city         string
	neighborhood string
	street       string
	service      string
	location     Location
}
