module v1

pub struct Ncm {
pub:
	codigo      string
	descricao   string
	data_inicio string
	data_fim    string
	tipo_ato    string
	numero_ato  string
	ano_ato     string
}
