module v1

// Quadro de Sócios e Administradores da empresa.
pub struct Qsa {
	pub:
	pais                                    string
	nome_socio                              string
	codigo_pais                             int
	faixa_etaria                            string
	cnpj_cpf_do_socio                       string
	qualificacao_socio                      string
	codigo_faixa_etaria                     int
	data_entrada_sociedade                  string
	identificador_de_socio                  int
	cpf_representante_legal                 string
	nome_representante_legal                string
	codigo_qualificacao_socio               int
	qualificacao_representante_legal        string
	codigo_qualificacao_representante_legal int
}
