module v1

pub struct Clima {
pub:
	data          string
	condicao      string
	min           int
	max           int
	indice_uv     int
	condicao_desc string
}
