module v1

import time

pub struct FeriadosNacional {
pub:
	date time.Time
	name string
	@type string
}
