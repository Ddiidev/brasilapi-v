module v2

pub struct Location {
	pub:
	@type       string
	coordinates Coordinates
}
