module v1

// Exemplo dos campos:<br/>
// codigo: Código da tabela de referência <br/>
// mes: Nome do mês/ano da tabela de referência<br/>
pub struct FipeTabelaReferencia {
pub:
	codigo int
	mes    string
}
